version https://git-lfs.github.com/spec/v1
oid sha256:893269fdccd2dc147e8570519f35308ac5e5460ad7f54bf673b3c31e9a8259de
size 2339
