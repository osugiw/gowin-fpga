version https://git-lfs.github.com/spec/v1
oid sha256:00d143e3b4226cb8ac7418bab35b9ea6f3a963e81fd0f2f7f3109844f4bde2c6
size 3219
