version https://git-lfs.github.com/spec/v1
oid sha256:39bfb925aa9600c0ce97a66fa28db792760a74fc1996999a2832de516649e033
size 1208
