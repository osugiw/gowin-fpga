version https://git-lfs.github.com/spec/v1
oid sha256:671d244e5a01dad9076059b777f1433ea6998442871f5f6fd72f28f2b40fe9b8
size 338
