version https://git-lfs.github.com/spec/v1
oid sha256:1e45e87703e2ab1790c13235822e8889fb016ad4c11cd9e5def0980d26a24637
size 4908
