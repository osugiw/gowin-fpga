version https://git-lfs.github.com/spec/v1
oid sha256:0e3a35ccb3e934eecfcd3916c5dac9ef269abea21472d66ebd2660a9d25e6a13
size 4612
