version https://git-lfs.github.com/spec/v1
oid sha256:b55c3af4cfbbdb7bb0445d0ef4afc9477d80a108e3740bc847edbcb18a7b4c0e
size 15431
