version https://git-lfs.github.com/spec/v1
oid sha256:dedd552fa988d9e2875bdadc54f3c08d5041d54637da1ff565d46078eeb2ea89
size 2395
