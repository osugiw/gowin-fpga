version https://git-lfs.github.com/spec/v1
oid sha256:6c3e87c8221a5756393bdbff0c48988f03e4917e0f088b7cba5cda8d6e83f3ad
size 7753
