version https://git-lfs.github.com/spec/v1
oid sha256:b21ce083bcec51f21f8dd25dc3bbcc3cc302982b603d005e1e576fd70f7c353e
size 10015
