version https://git-lfs.github.com/spec/v1
oid sha256:06db25636caa6512f1013837f8173ea059bd97340fdaf8f32856d518e51cfe61
size 9015
