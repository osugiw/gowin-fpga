version https://git-lfs.github.com/spec/v1
oid sha256:0309686e03ad33b26c1fe4e0210e67f8d3025baa8424a86834b72f9066039e9a
size 4074
