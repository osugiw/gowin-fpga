version https://git-lfs.github.com/spec/v1
oid sha256:c151e2675ad97ef36254044e42657f2d758512d305040137859f9b8806135f64
size 4906
