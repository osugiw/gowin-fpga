version https://git-lfs.github.com/spec/v1
oid sha256:8f23b42acbb4f0bdb0ee0745ac9aea42d9e19267d50a476da9184bae6000bd24
size 2972
