version https://git-lfs.github.com/spec/v1
oid sha256:1c0616b883499f88acaa84638e0474227201cc1a2836e1eb2f110285c79ea7e7
size 13161
